module adder_it1_TB;

	// Inputs
	reg [31:0] op1;
	reg [31:0] op2;

	// Outputs
	wire [31:0] result;

	// Instantiate the Unit Under Test (UUT)
	adder_it1 uut (
		.op1(op1), 
		.op2(op2), 
		.result(result)
	);

	initial begin
		// Initialize Inputs
		op1 = 0; op2 = 0;
      #10;
		op1=32'b00111111101001100110011001100110;//1.3
		op2=32'b00111111100110011001100110011010;//1.2
       #10;
		op1=32'b00111111010000000000000000000000;//0.75
		op2=32'b01000000010100000000000000000000;//3.25
		#10;
		op1=32'b01000000100000111101011100001010;//4.12
		op2=32'b01000000011010011001100110011010;//3.65
		#10;
		op1=32'b01000001000010111000010100011111;//8.72
		op2=32'b01000000010011110101110000101001;//3.24
		#10;
		op1=32'b01000010111101100000000000000000;//123
		op2=32'b01000000101001101011100001010010;//5.21
	end
initial begin $monitor ("%0d: %b",$time,result);end
initial begin #220; $finish; end      
		
endmodule
//expected output-
//// 10:01000000001000000000000000000000
////20:01000000100000000000000000000000
////30:01000000111110001010001111010111
////40:01000001001111110101110000101001
////50:01000011000000000011010111000011
	

